module INVD1 ( I, ZN)
input I
output ZN

timing I ZN, 0.542299

module DFQD1 ( Q, CP, D)
input CP, D
output Q

timing CP Q, 4.8694715
timing D Q, 0.0

module FA1D1 (A, B, CI, S, CO)
input A,B,CI
output S,CO

timing A CO, 5.54625
timing B CO, 4.422249
timing CI CO, 2.3798745
timing A S, 5.1899495
timing B S, 4.788601
timing CI S, 2.366857

module AN2D1 (A1, A2, Z)
input A1, A2
output Z

timing A1 Z, 1.8132095
timing A2 Z, 1.910383

module HA1D1 (A,B,S,CO)
input A, B
output S, CO

timing A CO, 1.5263355
timing B CO, 1.6756295
timing A S, 2.4507395
timing B S, 1.8878555

module XOR2D0 (A1, A2, Z)
input A1, A2
output Z

timing A1 Z, 2.370939
timing A2 Z, 3.2775585

module OR2D0 (A1, A2, Z)
input A1, A2
output Z

timing A1 Z, 2.0793405
timing A2 Z, 2.2433725

module OAI21D0 (A1, A2, B, ZN)
input A1, A2, B
output ZN

timing A1 ZN, 1.3178325
timing A2 ZN, 1.445072
timing B ZN, 1.0256165

module NR2D0 (A1, A2, ZN)
input A1, A2
output ZN

timing A1 ZN, 1.098822
timing A2 ZN, 1.149696

module CKND2D0 (A1, A2, ZN)
input A1, A2
output ZN

timing A1 ZN, 0.8399025
timing A2 ZN, 0.902671

module CKND0 (I, ZN)
input I
output ZN

timing I ZN, 0.637329

module AN2D0 (A1, A2, Z)
input A1, A2
output Z

timing A1 Z, 1.7415265
timing A2 Z, 1.8459565

module AOI21D0 (A1, A2, B, ZN)
input A1, A2, B
output ZN

timing A1 ZN, 1.345285
timing A2 ZN, 1.5098155
timing B ZN, 1.3746805

module OA22D0 (A1, A2, B1, B2, Z)
input A1, A2, B1, B2
output Z

timing A1 Z, 2.541883
timing A2 Z, 2.678619
timing B1 Z, 3.0788745
timing B2 Z, 3.1133855

module AOI22D0 (A1, A2, B1, B2, ZN)
input A1, A2, B1, B2
output ZN

timing A1 ZN, 1.322851
timing A2 ZN, 1.413906
timing B1 ZN, 1.7134165
timing B2 ZN, 1.802058

module AO21D0 (A1, A2, B, Z)
input A1, A2, B	
output Z

timing A1 Z, 2.5068275
timing A2 Z, 2.696815
timing B Z, 2.373018

module MUX2ND0 (I0, I1, S, ZN)
input I0, I1, S
output ZN

timing I0 ZN, 1.5642995
timing I1 ZN, 1.276669
timing S ZN, 2.072006

module AO22D0 (A1, A2, B1, B2, Z)
input A1, A2, B1, B2
output Z

timing A1 Z, 2.4386245
timing A2 Z, 2.6152235
timing B1 Z, 2.9511045
timing B2 Z, 3.0074175

module MAOI22D0 (A1, A2, B1, B2, ZN)
input A1, A2, B1, B2
output ZN

timing A1 ZN, 1.2523185
timing A2 ZN, 1.4282975
timing B1 ZN, 2.790838
timing B2 ZN, 2.921449

module OAI22D0 (A1, A2, B1, B2, ZN)
input A1, A2, B1, B2	
output ZN

timing A1 ZN, 1.4234735
timing A2 ZN, 1.492425
timing B1 ZN, 1.8116695
timing B2 ZN, 1.891133

module OA21D0 (A1, A2, B, Z)
input A1, A2, B
output Z

timing A1 Z, 2.507539
timing A2 Z, 2.646905
timing B Z, 1.9726225

module AOI22D1 (A1, A2, B1, B2, ZN)
input A1, A2, B1, B2
output ZN

timing A1 ZN, 1.322851
timing A2 ZN, 1.413906
timing B1 ZN, 1.7134165
timing B2 ZN, 1.802058

module XNR2D0 (A1, A2, ZN)
input A1, A2
output ZN

timing A1 ZN, 2.45697
timing A2 ZN, 3.307295

module MUX2D0 (I0, I1, S, Z)
input I0, I1, S
output Z

timing I0 Z, 3.0324515
timing I1 Z, 2.917908
timing S Z, 2.369111

module MOAI22D0 (A1, A2, B1, B2, ZN)
input A1, A2, B1, B2
output ZN

timing A1 ZN, 1.270133
timing A2 ZN, 1.4422855
timing B1 ZN, 2.1256305
timing B2 ZN, 2.2049545


module XOR4D1 (A1, A2, A3, A4, Z)
input A1, A2, A3, A4
output Z

timing A1 Z, 6.2737035
timing A2 Z, 6.539095
timing A3 Z, 6.488074
timing A4 Z, 5.9022865

module BUFFD1 (I, Z)
input I
output Z

timing I Z, 1.438696

module NR2D2 (A1, A2, ZN)
input A1, A2
output ZN

timing A1 ZN, 0.6748165
timing A2 ZN, 0.8203675

module BUFFD2 (I, Z)
input I
output Z

timing I Z, 1.2963915

module CKAN2D0 (A1, A2, Z)
input A1, A2
output Z

timing A1 Z, 1.8282275
timing A2 Z, 1.945969

module ND2D2 (A1, A2, ZN)
input A1, A2
output ZN

timing A1 ZN, 0.5640225
timing A2 ZN, 0.6667065

module OAI21D1 (A1, A2, B, ZN)
input A1, A2, B
output ZN

timing A1 ZN, 1.0190875
timing A2 ZN, 1.1698495
timing B ZN, 0.8797345

module ND2D1 (A1, A2, ZN)
input A1, A2
output ZN

timing A1 ZN, 0.7169115
timing A2 ZN, 0.7915985

module CKBD1 (I, Z)
input I
output Z

timing I Z, 1.2199855

module OR2D1 (A1, A2, Z)
input A1, A2
output Z

timing A1 Z, 1.8076425
timing A2 Z, 1.9552815

module CKND1 (I, ZN)
input I
output ZN

timing I ZN, 0.5560075

module INVD2 (I, ZN)
input I
output ZN

timing I ZN, 0.4735345

module AN2XD1 (A1, A2, Z)
input A1, A2
output Z

timing A1 Z, 1.466989
timing A2 Z, 1.584859

module NR2XD1 (A1, A2, ZN)
input A1, A2
output ZN

timing A1 ZN, 0.643466
timing A2 ZN, 0.8141785

module MUX4D1 (I0, I1, I2, I3, S0, S1, Z)
input I0, I1, I2, I3, S0, S1
output Z

timing I0 Z, 5.464088
timing I1 Z, 4.5712725
timing I2 Z, 5.7099275
timing I3 Z, 4.6643495
timing S0 Z, 4.7700715
timing S1 Z, 3.0733095

module INVD3 (I, ZN)
input I
output ZN

timing I ZN, 0.4568515

module AOI21D1 (A1, A2, B, ZN)
input A1, A2, B
output ZN

timing A1 ZN, 1.009721
timing A2 ZN, 1.1561905
timing B ZN, 1.0921565
