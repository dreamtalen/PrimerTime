
module c1355 ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, 
        G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, 
        G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, 
        G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, 
        G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
        G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, 
        G7, G8, G9 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200;

  XOR2D0 U127 ( .A1(n95), .A2(G32), .Z(G1355) );
  CKND2D0 U128 ( .A1(n96), .A2(n97), .ZN(n95) );
  XOR2D0 U129 ( .A1(n98), .A2(G31), .Z(G1354) );
  CKND2D0 U130 ( .A1(n96), .A2(n99), .ZN(n98) );
  XOR2D0 U131 ( .A1(n100), .A2(G30), .Z(G1353) );
  CKND2D0 U132 ( .A1(n96), .A2(n101), .ZN(n100) );
  XOR2D0 U133 ( .A1(n102), .A2(G29), .Z(G1352) );
  CKND2D0 U134 ( .A1(n96), .A2(n103), .ZN(n102) );
  AN2D0 U135 ( .A1(n104), .A2(n105), .Z(n96) );
  NR2D0 U136 ( .A1(n106), .A2(n107), .ZN(n104) );
  XOR2D0 U137 ( .A1(n108), .A2(G28), .Z(G1351) );
  CKND2D0 U138 ( .A1(n109), .A2(n97), .ZN(n108) );
  XOR2D0 U139 ( .A1(n110), .A2(G27), .Z(G1350) );
  CKND2D0 U140 ( .A1(n109), .A2(n99), .ZN(n110) );
  XOR2D0 U141 ( .A1(n111), .A2(G26), .Z(G1349) );
  CKND2D0 U142 ( .A1(n109), .A2(n101), .ZN(n111) );
  XOR2D0 U143 ( .A1(n112), .A2(G25), .Z(G1348) );
  CKND2D0 U144 ( .A1(n109), .A2(n103), .ZN(n112) );
  AN2D0 U145 ( .A1(n113), .A2(n114), .Z(n109) );
  NR2D0 U146 ( .A1(n115), .A2(n116), .ZN(n114) );
  CKND2D0 U147 ( .A1(n117), .A2(n118), .ZN(n116) );
  NR2D0 U148 ( .A1(n107), .A2(n119), .ZN(n113) );
  XNR2D0 U149 ( .A1(G24), .A2(n120), .ZN(G1347) );
  NR2D0 U150 ( .A1(n121), .A2(n122), .ZN(n120) );
  XNR2D0 U151 ( .A1(G23), .A2(n123), .ZN(G1346) );
  NR2D0 U152 ( .A1(n124), .A2(n122), .ZN(n123) );
  XNR2D0 U153 ( .A1(G22), .A2(n125), .ZN(G1345) );
  NR2D0 U154 ( .A1(n126), .A2(n122), .ZN(n125) );
  XNR2D0 U155 ( .A1(G21), .A2(n127), .ZN(G1344) );
  NR2D0 U156 ( .A1(n128), .A2(n122), .ZN(n127) );
  CKND2D0 U157 ( .A1(n129), .A2(n106), .ZN(n122) );
  AN2D0 U158 ( .A1(n107), .A2(n105), .Z(n129) );
  NR2D0 U159 ( .A1(n130), .A2(n115), .ZN(n105) );
  CKND2D0 U160 ( .A1(n119), .A2(n131), .ZN(n130) );
  XOR2D0 U161 ( .A1(n132), .A2(G20), .Z(G1343) );
  CKND2D0 U162 ( .A1(n133), .A2(n97), .ZN(n132) );
  XOR2D0 U163 ( .A1(n134), .A2(G19), .Z(G1342) );
  CKND2D0 U164 ( .A1(n133), .A2(n99), .ZN(n134) );
  XOR2D0 U165 ( .A1(n135), .A2(G18), .Z(G1341) );
  CKND2D0 U166 ( .A1(n133), .A2(n101), .ZN(n135) );
  XOR2D0 U167 ( .A1(n136), .A2(G17), .Z(G1340) );
  CKND2D0 U168 ( .A1(n133), .A2(n103), .ZN(n136) );
  AN2D0 U169 ( .A1(n137), .A2(n138), .Z(n133) );
  NR2D0 U170 ( .A1(n139), .A2(n131), .ZN(n138) );
  NR2D0 U171 ( .A1(n115), .A2(n140), .ZN(n137) );
  OAI21D0 U172 ( .A1(n121), .A2(n126), .B(n141), .ZN(n115) );
  AOI22D0 U173 ( .A1(n103), .A2(n142), .B1(n99), .B2(n143), .ZN(n141) );
  OR2D0 U174 ( .A1(n143), .A2(n99), .Z(n142) );
  XOR2D0 U175 ( .A1(n144), .A2(G16), .Z(G1339) );
  CKND2D0 U176 ( .A1(n145), .A2(n119), .ZN(n144) );
  XOR2D0 U177 ( .A1(n146), .A2(G15), .Z(G1338) );
  CKND2D0 U178 ( .A1(n145), .A2(n118), .ZN(n146) );
  XOR2D0 U179 ( .A1(n147), .A2(G14), .Z(G1337) );
  CKND2D0 U180 ( .A1(n145), .A2(n117), .ZN(n147) );
  XOR2D0 U181 ( .A1(n148), .A2(G13), .Z(G1336) );
  CKND2D0 U182 ( .A1(n145), .A2(n107), .ZN(n148) );
  AN2D0 U183 ( .A1(n149), .A2(n150), .Z(n145) );
  NR2D0 U184 ( .A1(n126), .A2(n103), .ZN(n149) );
  XOR2D0 U185 ( .A1(n151), .A2(G12), .Z(G1335) );
  CKND2D0 U186 ( .A1(n152), .A2(n119), .ZN(n151) );
  XOR2D0 U187 ( .A1(n153), .A2(G11), .Z(G1334) );
  CKND2D0 U188 ( .A1(n152), .A2(n118), .ZN(n153) );
  XOR2D0 U189 ( .A1(n154), .A2(G10), .Z(G1333) );
  CKND2D0 U190 ( .A1(n152), .A2(n117), .ZN(n154) );
  XOR2D0 U191 ( .A1(n155), .A2(G9), .Z(G1332) );
  CKND2D0 U192 ( .A1(n152), .A2(n107), .ZN(n155) );
  AN2D0 U193 ( .A1(n156), .A2(n157), .Z(n152) );
  NR2D0 U194 ( .A1(n97), .A2(n158), .ZN(n157) );
  CKND2D0 U195 ( .A1(n99), .A2(n101), .ZN(n158) );
  CKND0 U196 ( .I(n124), .ZN(n99) );
  NR2D0 U197 ( .A1(n159), .A2(n103), .ZN(n156) );
  CKND0 U198 ( .I(n128), .ZN(n103) );
  XOR2D0 U199 ( .A1(n160), .A2(G8), .Z(G1331) );
  CKND2D0 U200 ( .A1(n161), .A2(n119), .ZN(n160) );
  XOR2D0 U201 ( .A1(n162), .A2(G7), .Z(G1330) );
  CKND2D0 U202 ( .A1(n161), .A2(n118), .ZN(n162) );
  XOR2D0 U203 ( .A1(n163), .A2(G6), .Z(G1329) );
  CKND2D0 U204 ( .A1(n161), .A2(n117), .ZN(n163) );
  XOR2D0 U205 ( .A1(n164), .A2(G5), .Z(G1328) );
  CKND2D0 U206 ( .A1(n161), .A2(n107), .ZN(n164) );
  AN2D0 U207 ( .A1(n165), .A2(n150), .Z(n161) );
  NR2D0 U208 ( .A1(n166), .A2(n159), .ZN(n150) );
  CKND2D0 U209 ( .A1(n97), .A2(n124), .ZN(n166) );
  CKND0 U210 ( .I(n121), .ZN(n97) );
  NR2D0 U211 ( .A1(n128), .A2(n101), .ZN(n165) );
  CKND0 U212 ( .I(n126), .ZN(n101) );
  XOR2D0 U213 ( .A1(n167), .A2(G4), .Z(G1327) );
  CKND2D0 U214 ( .A1(n168), .A2(n119), .ZN(n167) );
  CKND0 U215 ( .I(n169), .ZN(n119) );
  XOR2D0 U216 ( .A1(n170), .A2(G3), .Z(G1326) );
  CKND2D0 U217 ( .A1(n168), .A2(n118), .ZN(n170) );
  XOR2D0 U218 ( .A1(n171), .A2(G2), .Z(G1325) );
  CKND2D0 U219 ( .A1(n168), .A2(n117), .ZN(n171) );
  CKND0 U220 ( .I(n106), .ZN(n117) );
  XOR2D0 U221 ( .A1(n172), .A2(G1), .Z(G1324) );
  CKND2D0 U222 ( .A1(n168), .A2(n107), .ZN(n172) );
  AN2D0 U223 ( .A1(n173), .A2(n174), .Z(n168) );
  NR2D0 U224 ( .A1(n124), .A2(n128), .ZN(n174) );
  XOR4D1 U225 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .Z(n128) );
  XOR4D1 U226 ( .A1(G21), .A2(G17), .A3(G29), .A4(G25), .Z(n178) );
  CKND2D0 U227 ( .A1(G37), .A2(G41), .ZN(n177) );
  XOR4D1 U228 ( .A1(n179), .A2(n176), .A3(n180), .A4(n181), .Z(n124) );
  XOR4D1 U229 ( .A1(G23), .A2(G19), .A3(G31), .A4(G27), .Z(n181) );
  CKND2D0 U230 ( .A1(G39), .A2(G41), .ZN(n180) );
  XOR4D1 U231 ( .A1(G4), .A2(G3), .A3(G1), .A4(G2), .Z(n176) );
  NR2D0 U232 ( .A1(n143), .A2(n159), .ZN(n173) );
  OAI21D0 U233 ( .A1(n169), .A2(n106), .B(n182), .ZN(n159) );
  AOI22D0 U234 ( .A1(n107), .A2(n183), .B1(n118), .B2(n140), .ZN(n182) );
  OR2D0 U235 ( .A1(n140), .A2(n118), .Z(n183) );
  CKND0 U236 ( .I(n131), .ZN(n118) );
  XOR4D1 U237 ( .A1(n184), .A2(n185), .A3(n186), .A4(n187), .Z(n131) );
  XOR4D1 U238 ( .A1(G15), .A2(G11), .A3(G7), .A4(G3), .Z(n187) );
  CKND2D0 U239 ( .A1(G35), .A2(G41), .ZN(n186) );
  CKND2D0 U240 ( .A1(n106), .A2(n169), .ZN(n140) );
  CKND0 U241 ( .I(n139), .ZN(n107) );
  XOR4D1 U242 ( .A1(n188), .A2(n185), .A3(n189), .A4(n190), .Z(n139) );
  XOR4D1 U243 ( .A1(G13), .A2(G1), .A3(G9), .A4(G5), .Z(n190) );
  CKND2D0 U244 ( .A1(G33), .A2(G41), .ZN(n189) );
  XOR4D1 U245 ( .A1(G20), .A2(G19), .A3(G17), .A4(G18), .Z(n185) );
  XOR4D1 U246 ( .A1(n191), .A2(n184), .A3(n192), .A4(n193), .Z(n106) );
  XOR4D1 U247 ( .A1(G14), .A2(G10), .A3(G6), .A4(G2), .Z(n193) );
  CKND2D0 U248 ( .A1(G34), .A2(G41), .ZN(n192) );
  XOR4D1 U249 ( .A1(G28), .A2(G27), .A3(G25), .A4(G26), .Z(n184) );
  XOR4D1 U250 ( .A1(n191), .A2(n188), .A3(n194), .A4(n195), .Z(n169) );
  XOR4D1 U251 ( .A1(G16), .A2(G12), .A3(G8), .A4(G4), .Z(n195) );
  CKND2D0 U252 ( .A1(G36), .A2(G41), .ZN(n194) );
  XOR4D1 U253 ( .A1(G24), .A2(G23), .A3(G21), .A4(G22), .Z(n188) );
  XOR4D1 U254 ( .A1(G32), .A2(G31), .A3(G29), .A4(G30), .Z(n191) );
  CKND2D0 U255 ( .A1(n121), .A2(n126), .ZN(n143) );
  XOR4D1 U256 ( .A1(n196), .A2(n179), .A3(n197), .A4(n198), .Z(n126) );
  XOR4D1 U257 ( .A1(G22), .A2(G18), .A3(G30), .A4(G26), .Z(n198) );
  CKND2D0 U258 ( .A1(G38), .A2(G41), .ZN(n197) );
  XOR4D1 U259 ( .A1(G9), .A2(G12), .A3(G10), .A4(G11), .Z(n179) );
  XOR4D1 U260 ( .A1(n196), .A2(n175), .A3(n199), .A4(n200), .Z(n121) );
  XOR4D1 U261 ( .A1(G24), .A2(G20), .A3(G32), .A4(G28), .Z(n200) );
  CKND2D0 U262 ( .A1(G41), .A2(G40), .ZN(n199) );
  XOR4D1 U263 ( .A1(G8), .A2(G7), .A3(G5), .A4(G6), .Z(n175) );
  XOR4D1 U264 ( .A1(G16), .A2(G15), .A3(G13), .A4(G14), .Z(n196) );
endmodule

